`include "defines.v"

module if_stage (
    input 	wire 					cpu_clk_50M,
    input 	wire 					cpu_rst_n,
    
    input   wire [ 1: 0         ]  jtsel,
    input   wire [`REG_BUS      ]  addr1,
    input   wire [`REG_BUS      ]  addr2,
    input   wire [`REG_BUS      ]  addr3,
    
    input   wire [`STALL_BUS    ]  stall,
    
    output  reg                    ice,
    output 	reg  [`INST_ADDR_BUS] 	pc,
    output 	wire [`INST_ADDR_BUS]	iaddr
    );
    
    wire [`INST_ADDR_BUS] pc_next; 
    assign pc_next = pc + 4;                  // ������һ��ָ��ĵ�ַ
    always @(*) begin
		if (cpu_rst_n == `RST_ENABLE || (stall[0] == `STOP && stall[1] == `NOSTOP)) begin
			ice <= `CHIP_DISABLE;		      // ��λ��ʱ��ָ��洢������  
		end else begin
			ice <= `CHIP_ENABLE; 		      // ��λ������ָ��洢��ʹ��
		end
	end

    always @(posedge cpu_clk_50M) begin
        if (cpu_rst_n == `RST_ENABLE)
            pc <= `PC_INIT;                   // ָ��洢�����õ�ʱ��PC���ֳ�ʼֵ��MiniMIPS32������Ϊ0x00000000��
        else if (stall[0] == `NOSTOP) begin
            case (jtsel)
                2'b00: pc <= pc_next;
                2'b01: pc <= addr3;
                2'b10: pc <= addr1;
                2'b11: pc <= addr2;
                default: pc <= pc_next; // ָ��洢��ʹ�ܺ�PCֵÿʱ�����ڼ�4 
            endcase	
        end
    end
    
    assign iaddr = (ice == `CHIP_DISABLE) ? `PC_INIT :
                   (stall[0] == `STOP && stall[1] == `STOP) ? pc - 4 : pc;    // ��÷���ָ��洢���ĵ�ַ

endmodule